module Ssegtobin (Ssegnum1, Ssegnum2, signo1, operador, num1, num2, sig1, oper);
	input [20:0] Ssegnum1;
	input [20:0] Ssegnum2;
	input [6:0] signo1;
	input [6:0] operador;
	output [9:0] num1;
	output [9:0] num2;
	output  sig1;
	output  oper;
	
endmodule
